module gen_data(
    output [127:0] row0,
    output [127:0] row1
);

    assign row0 = " Happy New Year ";
    assign row1 = "      2025      ";

endmodule
